AXILiteSimRecipe/reset-storm.AXILiteSimRecipe.bsv