package IOCapAxi;

import IOCapAxi_Types :: *;
import IOCapAxi_Flits :: *;
import IOCapAxi_Exposers :: *;
import IOCapAxi_Checker3s :: *;
import IOCapAxi_KeyManagers :: *;
import IOCapAxi_KeyManager2s :: *;
import IOCapAxi_Windows :: *;
import IOCapAxi_Konata :: *; // Purely for KONATA_OFF

export IOCapAxi_Types :: *;
export IOCapAxi_Flits :: *;
export IOCapAxi_Exposers :: *;
export IOCapAxi_Checker3s :: *;
export IOCapAxi_KeyManagers :: *;
export IOCapAxi_KeyManager2s :: *;
export IOCapAxi_Windows :: *;
export IOCapAxi_Konata :: *;

endpackage